module xorg(output Y,input A, B); 
  xor(Y,A,B);
endmodule
