// Code your design here
module xnorg(output Y, input A, B);
    xnor(Y, A, B); 
endmodule
