
module notg(output Y, input A, B);
    not(Y, A, B); 
endmodule
