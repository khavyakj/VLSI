module andg(output Y,input A, B); 
  and(Y,A,B);
endmodule
