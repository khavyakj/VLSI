// Code your design here
module norg(output Y,input A, B); 
  nor(Y,A,B);
endmodule
